`default_nettype none

module decode(
    input  wire [79:0]  data,
    input  wire [4:0]   data_valid,
    output wire [191:0] instruction,
    output wire         instruction_valid
);



endmodule